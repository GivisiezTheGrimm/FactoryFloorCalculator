INFO:HDLCompiler:1061 - Parsing VHDL file "D:/FactoryFloorCalculator2025/vardisp.vhdl" into library work
INFO:ProjectMgmt - Parsing design hierarchy completed successfully.
